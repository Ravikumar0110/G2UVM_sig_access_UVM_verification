package pkg;
      import uvm_pkg::*;
   `include "uvm_macros.svh"
	
	`include "G2U_sig_access_transection.sv"
	`include "G2U_sig_access_sequence.sv"
	`include "G2U_sig_access_sequncer.sv"
	`include "G2U_sig_access_monitor.sv"
	`include "G2U_sig_access_driver.sv"
	`include "G2U_sig_access_agent.sv"
	`include "G2U_sig_access_scoreboard.sv"
	
    `include "G2U_sig_access_env.sv"
    `include "G2U_sig_access_test.sv"
  
endpackage